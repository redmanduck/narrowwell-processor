module forwarding_unit(
	forwarding_unit_if.haswell fwif
);

	always_comb: begin
		
	end

endmodule
