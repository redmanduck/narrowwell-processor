`ifndef FWD_IF_VH
`define FWD_IF_VH
`include "cpu_types_pkg.vh"

interface forwarding_unit_if;
  modport haswell(
    
  );
endinterface
`endif